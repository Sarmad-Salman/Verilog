module fa3b_t();
reg [2:0]a,b;
reg ci;
wire [2:0]s;
wire c;
fa3b fa3b1(s,c,a,b,ci);
initial
begin
#100; a[0]=0; a[1]=0; a[2]=0; b[0]=0; b[1]=0; b[2]=0; ci=0; 
#100; a[0]=0; a[1]=0; a[2]=1; b[0]=0; b[1]=0; b[2]=1; ci=0; 
#100; a[0]=0; a[1]=1; a[2]=0; b[0]=0; b[1]=1; b[2]=0; ci=0; 
#100; a[0]=0; a[1]=1; a[2]=1; b[0]=0; b[1]=1; b[2]=1; ci=0; 
#100; a[0]=1; a[1]=0; a[2]=0; b[0]=1; b[1]=0; b[2]=0; ci=0; 
#100; a[0]=1; a[1]=0; a[2]=1; b[0]=1; b[1]=0; b[2]=1; ci=0; 
#100; a[0]=1; a[1]=1; a[2]=0; b[0]=1; b[1]=1; b[2]=0; ci=0; 
#100; a[0]=1; a[1]=1; a[2]=1; b[0]=1; b[1]=1; b[2]=1; ci=0;
#100; a[0]=0; a[1]=0; a[2]=0; b[0]=0; b[1]=0; b[2]=0; ci=1; 
#100; a[0]=0; a[1]=0; a[2]=1; b[0]=0; b[1]=0; b[2]=1; ci=1; 
#100; a[0]=0; a[1]=1; a[2]=0; b[0]=0; b[1]=1; b[2]=0; ci=1; 
#100; a[0]=0; a[1]=1; a[2]=1; b[0]=0; b[1]=1; b[2]=1; ci=1; 
#100; a[0]=1; a[1]=0; a[2]=0; b[0]=1; b[1]=0; b[2]=0; ci=1; 
#100; a[0]=1; a[1]=0; a[2]=1; b[0]=1; b[1]=0; b[2]=1; ci=1; 
#100; a[0]=1; a[1]=1; a[2]=0; b[0]=1; b[1]=1; b[2]=0; ci=1; 
#100; a[0]=1; a[1]=1; a[2]=1; b[0]=1; b[1]=1; b[2]=1; ci=1;
end
endmodule